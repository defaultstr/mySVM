1 16.0 0.537667 0.888396
-1 16.0 0.910936 0.852047
1 0.756724011028752 -2.258847 -1.06887
1 0.8473544577976894 0.862173 -0.809499
-1 0.9461178552814278 3.10061 4.585491
1 0.8188222598038266 0.318765 -2.944284
-1 15.909776316756076 3.544212 1.333109
1 0.5940891482466459 -1.307688 1.43838
-1 6.620082756430406 1.257698 0.066977
1 16.0 3.578397 1.370299
-1 13.12209360801537 0.938418 1.561034
1 0.08911515174039779 2.769437 -1.711516
1 0.46736482429200915 -1.349887 -0.102242
1 8.590245978617281 3.034923 -0.241447
1 10.519464301621055 0.725404 0.319207
-1 1.259074594786511 0.597731 1.399673
-1 0.5270345313646614 0.577624 2.489965
1 16.0 1.489698 0.627707
1 4.582966779509721 1.409034 1.093266
-1 0.6806719202618255 1.822625 3.711888
-1 2.8946336338973957 1.803947 1.805876
-1 7.896172658587894 3.41931 -0.138355
-1 4.404420962813946 2.291584 1.160411
1 1.9262437651082045 1.630235 -1.113501
-1 0.2628364676729952 1.195534 2.960954
1 16.0 1.034693 1.53263
-1 0.618563336307521 2.835088 3.436697
-1 6.0509120355895485 1.756285 0.0391
-1 16.0 0.834156 0.792155
