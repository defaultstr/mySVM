1 16.0 2.475425 0.145701
-1 15.999999999999998 1.682104 -0.131938
1 16.0 0.518601 1.83153
-1 16.0 1.530073 0.648679
1 16.0 1.50699 0.716744
1 16.0 1.819261 -0.328955
-1 10.454063868199011 1.234679 0.137025
1 15.999999999999998 1.936217 0.164361
-1 16.0 0.443422 1.145362
1 16.0 -0.186022 2.3165
1 16.0 0.672957 0.657131
1 16.0 0.558986 0.967816
-1 16.0 0.012469 2.177779
-1 16.0 1.242448 0.441327
-1 16.0 1.603946 0.327512
1 16.0 1.574942 0.956892
1 16.0 -0.021959 1.591326
-1 16.0 -0.372809 1.858593
1 16.0 0.881268 1.46838
-1 16.0 2.023691 0.10336
-1 16.0 2.229446 0.113597
1 16.0 0.478973 1.567996
1 2.7806524842842424 2.300486 0.395484
1 16.0 1.013038 -0.193494
-1 16.0 0.911127 2.424461
-1 16.0 0.594584 0.959401
-1 16.0 1.250251 0.428623
-1 16.0 0.239763 1.877865
1 7.673411383914783 1.383134 1.310189
