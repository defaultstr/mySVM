1 16.0 0.537667 0.888396
-1 16.0 0.910936 0.852047
1 0.7561320816164634 -2.258847 -1.06887
1 0.8443086320893229 0.862173 -0.809499
-1 0.9453713711439202 3.10061 4.585491
1 0.8189649756413134 0.318765 -2.944284
-1 15.910321086869931 3.544212 1.333109
1 0.5941217421732619 -1.307688 1.43838
-1 6.602133087771384 1.257698 0.066977
1 16.0 3.578397 1.370299
-1 13.133213978081656 0.938418 1.561034
1 0.08885662937326035 2.769437 -1.711516
1 0.4673917262716759 -1.349887 -0.102242
1 8.591140339519557 3.034923 -0.241447
1 10.507654571177463 0.725404 0.319207
-1 1.2492866394817983 0.597731 1.399673
-1 0.5257286242837367 0.577624 2.489965
1 16.0 1.489698 0.627707
1 4.587193386413318 1.409034 1.093266
-1 0.679910810748116 1.822625 3.711888
-1 2.8942342245761825 1.803947 1.805876
-1 7.895391370572755 3.41931 -0.138355
-1 4.403183152244855 2.291584 1.160411
1 1.9278893428592283 1.630235 -1.113501
-1 0.26281170934020104 1.195534 2.960954
1 16.0 1.034693 1.53263
-1 0.6188493711924579 2.835088 3.436697
-1 6.063218000827868 1.756285 0.0391
-1 16.0 0.834156 0.792155
